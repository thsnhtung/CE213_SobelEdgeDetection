library verilog;
use verilog.vl_types.all;
entity Shift_Register_tb is
end Shift_Register_tb;
