library verilog;
use verilog.vl_types.all;
entity Loader_2_tb is
end Loader_2_tb;
