library verilog;
use verilog.vl_types.all;
entity Gradient_Loader_tb is
end Gradient_Loader_tb;
