library verilog;
use verilog.vl_types.all;
entity Gradient_tb is
end Gradient_tb;
