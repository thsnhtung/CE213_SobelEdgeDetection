library verilog;
use verilog.vl_types.all;
entity Add_row_column_1_tb is
end Add_row_column_1_tb;
