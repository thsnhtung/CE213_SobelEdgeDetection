library verilog;
use verilog.vl_types.all;
entity Sobel_tb is
end Sobel_tb;
