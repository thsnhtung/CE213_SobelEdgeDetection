library verilog;
use verilog.vl_types.all;
entity Loader_tb is
end Loader_tb;
