library verilog;
use verilog.vl_types.all;
entity convolu_tb is
end convolu_tb;
