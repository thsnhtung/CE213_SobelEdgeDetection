library verilog;
use verilog.vl_types.all;
entity Padding_tb is
end Padding_tb;
