library verilog;
use verilog.vl_types.all;
entity Controller is
    generic(
        S0              : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        S1              : vl_logic_vector(0 to 1) := (Hi0, Hi1);
        S2              : vl_logic_vector(0 to 1) := (Hi1, Hi0);
        S3              : vl_logic_vector(0 to 1) := (Hi1, Hi1)
    );
    port(
        \Begin\         : in     vl_logic;
        CLK             : in     vl_logic;
        Start           : in     vl_logic;
        isEnd           : in     vl_logic;
        Reset           : out    vl_logic;
        Enable          : out    vl_logic;
        Finish          : out    vl_logic;
        current_state   : out    vl_logic_vector(1 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of S0 : constant is 1;
    attribute mti_svvh_generic_type of S1 : constant is 1;
    attribute mti_svvh_generic_type of S2 : constant is 1;
    attribute mti_svvh_generic_type of S3 : constant is 1;
end Controller;
