library verilog;
use verilog.vl_types.all;
entity Fast_Fifo_tb is
end Fast_Fifo_tb;
