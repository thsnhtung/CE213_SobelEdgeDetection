library verilog;
use verilog.vl_types.all;
entity Register_tb is
end Register_tb;
